`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/27/2025 10:19:58 AM
// Design Name: 
// Module Name: Control_Unit_Top
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Control_Unit_Top(Op, RegWrite,ImmSrc, ALUSrc, MemWrite, ResultSrc, Branch, funct3, funct7, ALUControl);
input [6:0]Op, funct7;
input [2:0] funct3;
output RegWrite, ALUSrc, MemWrite, ResultSrc, Branch;
output [1:0]ImmSrc;
output [2:0]ALUControl;

wire [1:0]ALUOp;
Main_Decoder Main_Decoder(.Op(Op), .RegWrite(RegWrite), .ImmSrc(ImmSrc), .MemWrite(MemWrite), .ResultSrc(ResultSrc), .Branch(Branch), .ALUSrc(ALUSrc), .ALUOp(ALUOp));
ALU_Decoder ALU_Decoder(.ALUOp(ALUOp), .funct3(funct3), .funct7(funct7), .Op(Op), .ALUControl(ALUControl));

endmodule
